//`include "uvm_pkg.svh"

package rv_test_pkg;


//import uvm_pkg.sv
import uvm_pkg::*
  //`include "dp_interface.sv"
`include "uvm_macros.svh"
	//`include "uvm_macros.svh"
//`include "tb_defs.sv"
`include "rv_xtn.sv"
`include "rv_seq.sv"
`include "rv_sequencer.sv"
//`include "apb_agt_config.sv"
//`include "env_config.sv"
`include "rv_driver.sv"
`include "rv_monitor.sv"
`include "rv_agent.sv"


//`include "virtual_sequencer.sv"
//`include "virtual_seqs.sv"
`include "rv_sb.sv"

`include "rv_env.sv"
`include "rv_test.sv"
endpackage
